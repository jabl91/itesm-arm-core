----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:36:18 04/27/2012 
-- Design Name: 
-- Module Name:    rom_mod - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity rom_mod is
    Port ( addr : in  STD_LOGIC_VECTOR (6 downto 0);
           out_oc : out  STD_LOGIC_VECTOR (4 downto 0);
           out_dir : out  STD_LOGIC_VECTOR (6 downto 0);
           out_data : out  STD_LOGIC_VECTOR (3 downto 0)
			 );
end rom_mod;

architecture Behavioral of rom_mod is

signal rom_data : std_logic_vector(15 downto 0);
--Declaracion de un ROM de 128x16 bits
type romtable is array(0 to 127) of std_logic_vector(15 downto 0);

constant romdata : romtable := (


--	X"180A",X"181B",X"182C",X"183D",X"184E",X"185F",X"1909",X"0800",
--	X"0800",X"0800",X"0800",X"0800",X"0800",X"0800",X"0800",X"0800",	--15
--	X"0F05",X"0E00",X"01E0",X"0000",X"0000",X"0000",X"0000",X"0000", 	--23
--	X"0100",X"0600",X"0600",X"0600",X"0000",X"0000",X"0000",X"0800", 	--31
--	X"0800",X"0800",X"0300",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF"




	X"1701",X"0800",X"0800",X"0800",X"0800",X"0800",X"0800",X"0700",
	X"0700",X"1702",X"0A00",X"0B00",X"0C05",X"0D00",X"1000",X"1000",	--15
	X"0F05",X"0E00",X"01E0",X"0000",X"0000",X"0000",X"0000",X"0000", 	--23
	X"0100",X"0600",X"0600",X"0600",X"0000",X"0000",X"0000",X"0800", 	--31
	X"0800",X"0800",X"0300",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF"




--	X"1703",X"0800",X"1100",X"0A00",X"0600",X"0500",X"0000",X"0C00",
--	X"0D00",X"0E00",X"0F00",X"170A",X"0900",X"0A00",X"0B00",X"100F",
--	X"0700",X"1400",X"040A",X"22F0",X"1302",X"1301",X"1300",X"1601", --23
--	X"0100",X"0600",X"0600",X"0600",X"0000",X"0000",X"0000",X"0800", --31
--	X"0800",X"0800",X"0300",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",
--	X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"0000",X"FFFF"
	);


begin

	process(addr)
	begin
		rom_data <= romdata(to_integer(unsigned(addr)));
	end process;
	
	out_oc <= rom_data(12 downto 8);
	out_dir <=  rom_data(15 downto 13) & rom_data(7 downto 4);
	out_data <= rom_data(3 downto 0);

end Behavioral;

