--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:43:17 05/05/2012
-- Design Name:   
-- Module Name:   C:/Users/rage/Dropbox/Grupo de Trabajo/Procesador 4 bits/uP_4_bits/reg_a_tb.vhd
-- Project Name:  uP_4_bits
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: reg_a
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY reg_a_tb IS
END reg_a_tb;
 
ARCHITECTURE behavior OF reg_a_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT reg_a
    PORT(
         in_bus : INOUT  std_logic_vector(7 downto 0);
         in_ram : INOUT  std_logic_vector(7 downto 0);
         load_a : IN  std_logic;
         sel : IN  std_logic;
         clk : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal load_a : std_logic := '0';
   signal sel : std_logic := '0';
   signal clk : std_logic := '0';

	--BiDirs
   signal in_bus : std_logic_vector(7 downto 0);
   signal in_ram : std_logic_vector(7 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: reg_a PORT MAP (
          in_bus => in_bus,
          in_ram => in_ram,
          load_a => load_a,
          sel => sel,
          clk => clk
        );

    -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		in_bus <= "00000001";
		
		in_ram <= "11111000";

      wait for clk_period*10;
		
		load_a <= '1';
		
		wait for clk_period*2;
		
		load_a <= '0';
		
		sel <= '1';
		
		in_bus <= "00000100";

      -- insert stimulus here 

      wait;
   end process;

END;
